interface det_if (input bit clk);
    logic rstn;
    logic in;
    logic out;
endinterface //interfacename det_if (input bit clk);
